module top_module( 
    input a, 
    input b, 
    output out );
    
    and (out, a, b);

endmodule
